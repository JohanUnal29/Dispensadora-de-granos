`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:51:26 06/26/2023 
// Design Name: 
// Module Name:    Comparador_de_conteo 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

/*
 * Generated by Digital. Don't modify this file!
 * Any changes will be lost if this file is regenerated.
 */

module CompUnsigned #(
    parameter Bits = 1
)
(
    input [(Bits -1):0] a,
    input [(Bits -1):0] b,
    output \> ,
    output \= ,
    output \<
);
    assign \> = a > b;
    assign \= = a == b;
    assign \< = a < b;
endmodule


module Mux_2x1
(
    input [0:0] sel,
    input in_0,
    input in_1,
    output reg out
);
    always @ (*) begin
        case (sel)
            1'h0: out = in_0;
            1'h1: out = in_1;
            default:
                out = 'h0;
        endcase
    end
endmodule


module Comparador_de_conteo (
  input [3:0] Num_repeticiones,
  input X1,
  input [3:0] rise_count,
  output \Senal_frenado_maquina_estados 
);
  wire s0;
  CompUnsigned #(
    .Bits(4)
  )
  CompUnsigned_i0 (
    .a( Num_repeticiones ),
    .b( rise_count ),
    .\= ( s0 )
  );
  Mux_2x1 Mux_2x1_i1 (
    .sel( s0 ),
    .in_0( X1 ),
    .in_1( 1'b0 ),
    .out( \Se�al_frenado_maquina_estados  )
  );
endmodule
